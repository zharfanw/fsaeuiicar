* /media/mzharfanw/ZhardiskFile/Zharfan's Document/Project Document/EVProjectFSAE2019/Documentation/ShutdownSystem.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Min 26 Mei 2019 05:45:20  WIB

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
K1  42 39 ? 3 34 ? 42 4 FINDER-41.52		
D1  42 4 D		
Q1  3 36 42 MPSA92		
R1  ? 36 R		
K2  35 39 ? 34 40 ? 35 4 FINDER-41.52		
D2  35 4 D		
Q2  3 28 35 MPSA92		
R6  ? 28 R		
K3  47 39 ? 40 32 ? 47 4 FINDER-41.52		
D3  47 4 D		
Q4  3 49 47 MPSA92		
Q3  47 ? 49 MPSA42		
Reset1  ? 39 Conn_01x02		
ShutdownSeries1  32 19 Conn_01x02		
XU1  ? 42 10 4 ? 9 ? ? OP07		
R2  3 10 R		
R3  10 4 R		
R4  3 9 R		
R5  9 4 R		
XU2  ? 35 1 4 ? 2 ? ? OP07		
R7  3 1 R		
R8  1 4 R		
R9  3 2 R		
R10  2 4 R		
XU3  ? 47 25 4 ? 26 ? ? OP07		
R11  3 25 R		
R12  25 4 R		
R13  3 26 R		
R14  26 4 R		
IMDIndicator1  9 4 Conn_01x02		
BMSIndicator1  2 4 Conn_01x02		
BSPDIndicator1  26 4 Conn_01x02		
K4  ? ? ? 19 4 FINDER-40.51		
K5  ? ? ? ? ? ? 19 4 FINDER-41.52		

.end
